** Profile: "Startup-tran"  [ D:\Git\ishero\circuit_simulation\pspiceTI\TPS40170\TPS40170_PSPICE_TRANS\tps40170-pspicefiles\startup\tran.sim ] 

** Creating circuit file "tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../tps40170.lib" 
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\17.4.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1.8m 0 20n 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.OPTIONS ABSTOL= 10n
.OPTIONS ITL1= 1500
.OPTIONS ITL2= 400
.OPTIONS ITL4= 400
.OPTIONS VNTOL= 10u
.PROBE64 V(alias(*)) I(alias(*)) 
.INC "..\Startup.net" 


.END
